'parameter test
v1 1 0 dc (a) ac 'b'
r1 1 2 "c"
r2 2 0 {d}
.param a=1 b=2 c=3 d=4
.param
.print op v(nodes)
.op
.end
