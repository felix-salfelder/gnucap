*oscillator, .159 Hz.
C1 1 0 1 ic=5
L1 1 0 1

C2 2 0 1
L2 2 0 1 ic=5

.width out=80
* .options initsc 1
.print tran v(1) v(2) iter(0)
.tran .1 100 0 uic trace rejected
*.tran
*.tran
*.tran .1 100 0
.status notime
.tran .1 100 0 uic trace rejected
.status notime
.end
