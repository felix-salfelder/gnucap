'parameter test
v1 1 0 dc (a) ac b
r1 1 2 {a+b}
r2 2 0 d
.list
.param a=1 b=2 c=3 d=4
.list
.param
.print op v(nodes)
.op
.print ac v(nodes)
.ac
.end
