'inductance check, no tolerance
.options method traponly
V1   1  0  dc 1 ac 1  pulse iv=0,pv=1,rise=1,fall=1
L3   1  2  1.
R4   2  0  1.
R5   1  3  1.
C6   3  0  1.
E1   4  0  3  0  1.
rspice 4 0 1g
G1   5  0  3  0  1.
Rg   5  0  1.
.op
.print ac vm(2) vm(3) vm(4) vm(5) vp(2) vp(3) vp(4) vp(5)
.ac dec 1 .1 1
.print tran v(2) v(3) v(4) v(5)
.tran 1 10 0
.list
.status notime
.end
