.title mos3 inverter

.width out=550
.options initsc 1
*.options method traponly

.model nmos nmos level=3 vto=0.7
.model pmos pmos level=3 vto=-0.7

Mp1 3 2 1 1 PMOS W=8e-6 L=600e-9 
Mn1 3 2 0 0 NMOS W=8e-6 L=600e-9 

Mp2 4 2 1 1 PMOS W=8e-6 L=600e-9 
Mn2 4 2 0 0 NMOS W=8e-6 L=600e-9 
R2  4 0 10k

Mp3 5 2 1 1 PMOS W=8e-6 L=600e-9 
Mn3 5 2 0 0 NMOS W=8e-6 L=600e-9 
C3  5 0 1p

Mp4 6 2 1 1 PMOS W=8e-6 L=600e-9 
R4  6 0 5.6k

Mn5 7 2 0 0 NMOS W=8e-6 L=600e-9 
R5  7 1 5.6k

vdd 1 0 5
* vin 2 0 PWL (0 0, 1n 0, 3n 5, 10n 5, 12n 0, 20n 0)
vin 2 0 pulse iv=0 delay=1n rise=2n pv=5

.op

.print dc v(1) v(2) v(3) v(4) v(5) v(6) v(7)
.dc vin 0 5 .25

.print tran v(1) v(2) v(3) v(4) v(5) v(6) v(7) hidden(0) method(c*) dis(2)
+ method(Mp2.cg*) v(MP2.nodes)
.tran 0.1n 5n basic trace=a > bla.out
.tran 0.1n 5n basic trace=a

.status notime
.end
