'dctran test
V1   1  0  dc generator(1) ac 1
L3   1  2  dc 1. ac 1.
R4   2  0  dc 1. ac 1.
R5   1  3  dc 1. ac 1.
C6   3  0  dc 1. ac 1.
.options short=1p
.options initsc 1
.print tran iter(0)  v(nodes) control(0)
.tran 0 1 .1 trace rejected
.print ac v(nodes)
.ac .001 10 decade
.list
.status notime
.end
