'
V1  1  0  dc 1 ac 1
R1  1  2  10k
Yl1  2  0  100u
Vc2  3  0  1.
R2  1  4  10k
.vcg Rv2  4  0  3  0  100u
Vc3  5  0  2.
R3  1  6  5k
.vcg Rv3  6  0  5  0  100u
.print op v(2,3,4,5,6) iter(0)
.op trace iter
.delete Vc3
Vc3 5 0 sin freq=1k ampl=1 offset=1
.modify R3=10k
.print tran v(2,3,4,5,6) iter(0) control(0)
.tran 0 .001 .0001 trace iter
.status notime
.end
