# list

C1 0 1 5
C2 0 1 5 m=2
T1 0 1 2 3
T2 0 1 2 3 m=2
T3 0 1 2 3 z0=100 f=10meg
T4 0 1 2 3 z0=100 f=10meg m=2
.list
