'parameter test
v1 1 0 dc (a) ac b
r1 1 2 c
r2 2 0 c+1
.list
.param a=1 b=a+1 c=a+b d=c+1
.param
.print op v(nodes)
.op
.end
