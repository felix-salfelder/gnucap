spice

.subckt test na nb
r00 na n00 1
r01 na n01 1
r02 na n02 1
r03 na n03 1
r04 na n04 1
r05 na n05 1
r06 na n06 1
r07 na n07 1
r08 na n08 1
r09 na n09 1
r10 na n10 1
r12 na n12 1
r13 na n13 1
r14 na n14 1
r15 na n15 1
r16 na n16 1
r17 na n17 1
r18 na n18 1
r19 na n19 1
r20 na n20 1
r22 na n22 1
r23 na n23 1
r24 na n24 1
r25 na n25 1
r26 na n26 1
r27 na n27 1
r28 na n28 1
r29 na n29 1
r30 na n30 1
r32 na n32 1
r33 na n33 1
r34 na n34 1
r35 na n35 1
r36 na n36 1
r37 na n37 1
r38 na n38 1
r39 na n39 1
r40 na n40 1
r42 na n42 1
r43 na n43 1
r44 na n44 1
r45 na n45 1
r46 na n46 1
r47 na n47 1
r48 na n48 1
r49 na n49 1
r50 na n50 1
r52 na n52 1
r53 na n53 1
r54 na n54 1
r55 na n55 1
r56 na n56 1
r57 na n57 1
r58 na n58 1
r59 na n59 1
r60 na n60 1
r62 na n62 1
r63 na n63 1
r64 na n64 1
r65 na n65 1
r66 na n66 1
r67 na n67 1
r68 na n68 1
r69 na n69 1
r70 na n70 1
r72 na n72 1
r73 na n73 1
r74 na n74 1
r75 na n75 1
r76 na n76 1
r77 na n77 1
r78 na n78 1
r79 na n79 1
r80 na n80 1
r82 na n82 1
r83 na n83 1
r84 na n84 1
r85 na n85 1
r86 na n86 1
r87 na n87 1
r88 na n88 1
r89 na n89 1
r90 na n90 1
r92 na n92 1
r93 na n93 1
r94 na n94 1
r95 na n95 1
r96 na n96 1
r97 na n97 1
r98 na n98 1
r99 na n99 1

r100 na n100 1
r101 na n101 1
r102 na n102 1
r103 na n103 1
r104 na n104 1
r105 na n105 1
r106 na n106 1
r107 na n107 1
r108 na n108 1
r109 na n109 1
r110 na n110 1
r112 na n112 1
r113 na n113 1
r114 na n114 1
r115 na n115 1
r116 na n116 1
r117 na n117 1
r118 na n118 1
r119 na n119 1
r120 na n120 1
r122 na n122 1
r123 na n123 1
r124 na n124 1
r125 na n125 1
r126 na n126 1
r127 na n127 1
r128 na n128 1
r129 na n129 1
r130 na n130 1
r132 na n132 1
r133 na n133 1
r134 na n134 1
r135 na n135 1
r136 na n136 1
r137 na n137 1
r138 na n138 1
r139 na n139 1
r140 na n140 1
r142 na n142 1
r143 na n143 1
r144 na n144 1
r145 na n145 1
r146 na n146 1
r147 na n147 1
r148 na n148 1
r149 na n149 1
r150 na n150 1
r152 na n152 1
r153 na n153 1
r154 na n154 1
r155 na n155 1
r156 na n156 1
r157 na n157 1
r158 na n158 1
r159 na n159 1
r160 na n160 1
r162 na n162 1
r163 na n163 1
r164 na n164 1
r165 na n165 1
r166 na n166 1
r167 na n167 1
r168 na n168 1
r169 na n169 1
r170 na n170 1
r172 na n172 1
r173 na n173 1
r174 na n174 1
r175 na n175 1
r176 na n176 1
r177 na n177 1
r178 na n178 1
r179 na n179 1
r180 na n180 1
r182 na n182 1
r183 na n183 1
r184 na n184 1
r185 na n185 1
r186 na n186 1
r187 na n187 1
r188 na n188 1
r189 na n189 1
r190 na n190 1
r192 na n192 1
r193 na n193 1
r194 na n194 1
r195 na n195 1
r196 na n196 1
r197 na n197 1
r198 na n198 1
r199 na n199 1

c00 na n00 1
c01 na n01 1
c02 na n02 1
c03 na n03 1
c04 na n04 1
c05 na n05 1
c06 na n06 1
c07 na n07 1
c08 na n08 1
c09 na n09 1
c10 na n10 1
c12 na n12 1
c13 na n13 1
c14 na n14 1
c15 na n15 1
c16 na n16 1
c17 na n17 1
c18 na n18 1
c19 na n19 1
c20 na n20 1
c22 na n22 1
c23 na n23 1
c24 na n24 1
c25 na n25 1
c26 na n26 1
c27 na n27 1
c28 na n28 1
c29 na n29 1
c30 na n30 1
c32 na n32 1
c33 na n33 1
c34 na n34 1
c35 na n35 1
c36 na n36 1
c37 na n37 1
c38 na n38 1
c39 na n39 1
c40 na n40 1
c42 na n42 1
c43 na n43 1
c44 na n44 1
c45 na n45 1
c46 na n46 1
c47 na n47 1
c48 na n48 1
c49 na n49 1
c50 na n50 1
c52 na n52 1
c53 na n53 1
c54 na n54 1
c55 na n55 1
c56 na n56 1
c57 na n57 1
c58 na n58 1
c59 na n59 1
c60 na n60 1
c62 na n62 1
c63 na n63 1
c64 na n64 1
c65 na n65 1
c66 na n66 1
c67 na n67 1
c68 na n68 1
c69 na n69 1
c70 na n70 1
c72 na n72 1
c73 na n73 1
c74 na n74 1
c75 na n75 1
c76 na n76 1
c77 na n77 1
c78 na n78 1
c79 na n79 1
c80 na n80 1
c82 na n82 1
c83 na n83 1
c84 na n84 1
c85 na n85 1
c86 na n86 1
c87 na n87 1
c88 na n88 1
c89 na n89 1
c90 na n90 1
c92 na n92 1
c93 na n93 1
c94 na n94 1
c95 na n95 1
c96 na n96 1
c97 na n97 1
c98 na n98 1
c99 na n99 1
c100 na n100 1
c101 na n101 1
.ends

Xt 1 0 test
.list

.print op v(nodes) v(xT.nodes)
.print
.print op

.end
