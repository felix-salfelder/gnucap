spice

*.options trace
v1 n1 0 pulse iv=0 pv=1 rise=1m delay=1m width=3m fall=5m
v2 n3 0 pulse iv=0 pv=1 rise=1m delay=3m width=3m fall=5m

cd n1 n3 0

c1 n2 0 200n
r1 n1 n2 1k

c2 n4 0 200n
r2 n3 n4 1k

.list

.print tran v(nodes) method(c*) disc(nodes) hidden(0)
.options initsc 1
.tran 0 5m 5m basic trace=a

.stat notime

.echo traponly
.options method traponly
.options initsc -1
.tran 0 5m 5m trace=a

.stat notime
.end
